`default_nettype none
module top (
    // HW
    input clk, nrst,
    
    // Wrapper
    input cs,
    inout [33:0] gpio
);



endmodule