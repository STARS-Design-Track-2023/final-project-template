`default_nettype none
module tb_top (

);

endmodule